module ();
    input ;
    output ;

endmodule

