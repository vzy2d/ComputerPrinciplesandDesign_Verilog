module ();
input ;
output ;

endmodule

/*
-Notepad++自动补全-
module endmodule
assign wire reg
begin end
initial always
function endfunction
task endtask
case default endcase
parameter
posedge negedge
*/